// Copyright 2021 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_MIO_CLI_MACROS_SVH__
`define __UVMA_MIO_CLI_MACROS_SVH__





`endif // __UVMA_MIO_CLI_MACROS_SVH__
