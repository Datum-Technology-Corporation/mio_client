// Copyright 2021 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_MIO_CLI_ST_MACROS_SVH__
`define __UVME_MIO_CLI_ST_MACROS_SVH__





`endif // __UVME_MIO_CLI_ST_MACROS_SVH__
